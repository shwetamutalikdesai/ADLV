edftrtgvtr
